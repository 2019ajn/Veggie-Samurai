`timescale 1ns / 1ps
`default_nettype none

module katana_tracking(

);

endmodule

`default_nettype wire