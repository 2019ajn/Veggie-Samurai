`timescale 1ns / 1ps
`default_nettype none

module game_logic_tb(
	
	);

endmodule

`default_nettype wire