`timescale 1ns / 1ps
`default_nettype none

module parabolic (
    input wire clk_in, rst_in, split_in, veggie_gone_in,
    output logic[2:0] x_speed_out, y_speed_out,
    output logic up // what is this for again?
);


endmodule

`default_nettype wire